//----------------------------------//
// Breakout Files
// y-block.v
// David J. Morvay
// ECEN 4856
// Fall 2020
//----------------------------------//

module y_block(pix_x, pix_y, block_on);
input [10:0] pix_x, pix_y;
output block_on;
// Square Y
localparam BALL_SIZE = 64;
// Y left, right boundary
wire [10:0] y_x_l = 368;
wire [10:0] y_x_r = y_x_l + BALL_SIZE - 1;
// Y top, bottom boundary 
wire [10:0] y_y_t = 268; 
wire [10:0] y_y_b = y_y_t + BALL_SIZE - 1;

// Y
wire [5:0] rom_addr, rom_col;
reg [63:0] rom_data;
wire rom_bit;

// "Y" image ROM
always @*
case (rom_addr)
	6'h0: rom_data =   64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
	6'h1: rom_data =   64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;	
	6'h2: rom_data =   64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;
	6'h3: rom_data =   64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;
	6'h4: rom_data =   64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;	
	6'h5: rom_data =   64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;		
	6'h6: rom_data =   64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;		
	6'h7: rom_data =   64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;	 
	6'h8: rom_data =   64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;
	6'h9: rom_data =   64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;
	6'hA: rom_data =   64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;	
	6'hB: rom_data =   64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;		
	6'hC: rom_data =   64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;		
	6'hD: rom_data =   64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;	 
	6'hE: rom_data =   64'b11001111_11111111_11111111_11110000_11111111_11111111_11111111_11110011; 
	6'hF: rom_data =   64'b11001111_11111111_11111111_11110000_11111111_11111111_11111111_11110011;
	6'h10: rom_data =  64'b11001111_11111111_11111111_11110000_11111111_11111111_11111111_11110011;
	6'h11: rom_data =  64'b11001111_11111111_11111111_11110000_11111111_11111111_11111111_11110011;
	6'h12: rom_data =  64'b11001111_11111111_11111111_11110000_11111111_11111111_11111111_11110011; 
	6'h13: rom_data =  64'b11001111_11111111_11111111_11110000_11111111_11111111_11111111_11110011;
	6'h14: rom_data =  64'b11001111_11111111_11111111_11110000_11111111_11111111_11111111_11110011;
	6'h15: rom_data =  64'b11001111_11111111_11111111_11110000_11111111_11111111_11111111_11110011;
	6'h16: rom_data =  64'b11000000_00111111_11111111_00000000_00000011_11111111_11111100_00000011;
	6'h17: rom_data =  64'b11000000_00011111_11111111_10000000_00000111_11111111_11111000_00000011;
	6'h18: rom_data =  64'b11000000_00001111_11111111_11000000_00001111_11111111_11110000_00000011; 
	6'h19: rom_data =  64'b11000000_00000111_11111111_11100000_00011111_11111111_11100000_00000011;
	6'h1A: rom_data =  64'b11000000_00000011_11111111_11110000_00111111_11111111_11000000_00000011;
	6'h1B: rom_data =  64'b11000000_00000001_11111111_11111000_01111111_11111111_10000000_00000011;
	6'h1C: rom_data =  64'b11000000_00000000_11111111_11111100_11111111_11111111_00000000_00000011;
	6'h1D: rom_data =  64'b11000000_00000000_01111111_11111111_11111111_11111110_00000000_00000011;	
	6'h1E: rom_data =  64'b11000000_00000000_00111111_11111111_11111111_11111100_00000000_00000011;
	6'h1F: rom_data =  64'b11000000_00000000_00011111_11111111_11111111_11111000_00000000_00000011;	
	6'h20: rom_data =  64'b11000000_00000000_00001111_11111111_11111111_11110000_00000000_00000011;	
	6'h21: rom_data =  64'b11000000_00000000_00000111_11111111_11111111_11100000_00000000_00000011;	
	6'h22: rom_data =  64'b11000000_00000000_00000011_11111111_11111111_11000000_00000000_00000011;	
	6'h23: rom_data =  64'b11000000_00000000_00000001_11111111_11111111_10000000_00000000_00000011;
	6'h24: rom_data =  64'b11000000_00000000_00000000_11111111_11111111_00000000_00000000_00000011;			
	6'h25: rom_data =  64'b11000000_00000000_00000000_01111111_11111110_00000000_00000000_00000011;
	6'h26: rom_data =  64'b11000000_00000000_00000000_00111111_11111100_00000000_00000000_00000011;
	6'h27: rom_data =  64'b11000000_00000000_00000000_00111111_11111100_00000000_00000000_00000011;
	6'h28: rom_data =  64'b11000000_00000000_00000000_00111111_11111100_00000000_00000000_00000011;
	6'h29: rom_data =  64'b11000000_00000000_00000000_00111111_11111100_00000000_00000000_00000011;
	6'h2A: rom_data =  64'b11000000_00000000_00000000_00111111_11111100_00000000_00000000_00000011; 
	6'h2B: rom_data =  64'b11000000_00000000_00000000_00111111_11111100_00000000_00000000_00000011; 
	6'h2C: rom_data =  64'b11000000_00000000_00111111_11111111_11111111_11111100_00000000_00000011;
	6'h2D: rom_data =  64'b11000000_00000000_00111111_11111111_11111111_11111100_00000000_00000011;
	6'h2E: rom_data =  64'b11000000_00000000_00111111_11111111_11111111_11111100_00000000_00000011;
	6'h2F: rom_data =  64'b11000000_00000000_00111111_11111111_11111111_11111100_00000000_00000011;
	6'h30: rom_data =  64'b11000000_00000000_00111111_11111111_11111111_11111100_00000000_00000011;
	6'h31: rom_data =  64'b11000000_00000000_00111111_11111111_11111111_11111100_00000000_00000011;
	6'h32: rom_data =  64'b11000000_00000000_00111111_11111111_11111111_11111100_00000000_00000011;
	6'h33: rom_data =  64'b11000000_00000000_00111111_11111111_11111111_11111100_00000000_00000011;
	6'h34: rom_data =  64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;	
	6'h35: rom_data =  64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;
	6'h36: rom_data =  64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;
	6'h37: rom_data =  64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;
	6'h38: rom_data =  64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;
	6'h39: rom_data =  64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;
	6'h3A: rom_data =  64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;
	6'h3B: rom_data =  64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;
	6'h3C: rom_data =  64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;
	6'h3D: rom_data =  64'b11000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;
	6'h3E: rom_data =  64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
	6'h3F: rom_data =  64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;		

	
	//   ****************************************************************
	//   ****************************************************************
	//   **                                                            **
	//   **                                                            **
	//   **                                                            **
	//   **                                                            **
	//   **                                                            **
	//   **                                                            **
	//   **                                                            **
	//   **                                                            **
	//   **                                                            **
	//   **                                                            **
	//   **                                                            **
	//   **                                                            **
	//   **  ************************    ****************************  **
	//   **  ************************    ****************************  **
	//   **  ************************    ****************************  **
	//   **  ************************    ****************************  **
	//   **  ************************    ****************************  **
	//   **  ************************    ****************************  **
	//   **  ************************    ****************************  **
	//   **  ************************    ****************************  **
	//   **        **************              ****************        **
	//   **         **************            ****************         **
	//   **          **************          ****************          **
	//   **           **************        ****************           **
	//   **            **************      ****************            **	
	//   **             **************    ****************             **
	//   **              **************  ****************              **
	//   **               ******************************               **
	//   **                ****************************                **
	//   **                 **************************                 **
	//   **                  ************************                  **
	//   **                   **********************                   **	
	//   **                    ********************                    **
	//   **                     ******************                     **
	//   **                      ****************                      **
	//   **                       **************                       **
	//   **                        ************                        **
	//   **                        ************                        **
	//   **                        ************                        **
	//   **                        ************                        **
	//   **                        ************                        **
	//   **                        ************                        **
	//   **                ****************************                **
	//   **                ****************************                **
	//   **                ****************************                **
	//   **                ****************************                **
	//   **                ****************************                **
	//   **                ****************************                **
	//   **                ****************************                **
	//   **                ****************************                **	
	//   **                                                            **
	//   **                                                            **
	//   **                                                            **
	//   **                                                            **
	//   **                                                            **
	//   **                                                            **
	//   **                                                            **
	//   **                                                            **
	//   **                                                            **
	//   **                                                            **
	//   ****************************************************************
	//   ****************************************************************
					
endcase

//---------------------------- Ball Body --------------------------------------------------//

// Pixel within square box
assign sq_y_on = (y_x_l <= pix_x) && (pix_x <= y_x_r) && (y_y_t <= pix_y) && (pix_y <= y_y_b);
// Map current pixel location to ROM addr/col
assign rom_addr = pix_y[5:0] - y_y_t[5:0];
assign rom_col = pix_x[5:0] - y_x_l[5:0];
assign rom_bit = rom_data[rom_col];
// Pixel within "Y"
assign block_on = sq_y_on && rom_bit;

endmodule
